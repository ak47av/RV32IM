`timescale 1ns / 1ps

module SSplitter(
    input  logic [31:0] ins,
    output logic [6:0] opcode,
    output logic  [4:0] imm4_0,
    output logic  [2:0] funct3,
    output logic  [4:0] rs1,
    output logic  [4:0] rs2,
    output logic  [6:0] imm11_5
    );
    
    assign {imm11_5, rs2, rs1, funct3, imm4_0, opcode} = ins;
    
endmodule
